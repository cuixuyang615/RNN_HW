`ifndef ALU_defines
`define ALU_defines

`define ALUADD      4'd0
`define ALUSUB      4'd1
`define ALUAND      4'd2
`define ALUOR       4'd3
`define ALUMUL      4'd4
`define ALUSLT      4'd5      //could use sub to determine? //`define ALUDIV      4'd5
`define ALUFADD     4'd6
`define ALUFSUB     4'd7
`define ALUFMUL     4'd8
`define ALUFDIV     4'd9      //disabled
`define ALUFADDM    4'd10
`define ALUFDOTM    4'd11
`define ALUFSUMM    4'd12
`define ALUFSIGM    4'd13
`define ALUFTANHM   4'd14
`define ALUINVALID  4'd15



`endif 
